package alu_type is

    -- ALU OP Type
    type alu_op_t is (
        ALU_ADD,
        ALU_SUB
    );

end alu_type;
